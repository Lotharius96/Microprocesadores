-- File Name   : lfsr_pkg.vhd
------------------------------------------------------------------
library ieee;
    use ieee.std_logic_1164.all;
    use ieee.std_logic_textio.all;
	 use ieee.numeric_std.ALL;
    use std.textio.all;
    
package lfsr_pkg is
	
    constant LFSR_W : natural := 6;		-- LFSR width
	
end lfsr_pkg; 
